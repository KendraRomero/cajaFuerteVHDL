library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity SIETE_SEGMENTOS is port(
	ENTRADA : in std_logic_vector(3 downto 0);
	SALIDA_SIETE_SEGMENTOS : out std_logic_vector(6 downto 0)
); end SIETE_SEGMENTOS;

architecture LOGICA_SIETE_SEGMENTOS of SIETE_SEGMENTOS is

begin
	with ENTRADA select SALIDA_SIETE_SEGMENTOS <=
		"1000000" when "0000",
		"1111001" when "0001",
		"0100100" when "0010",
		"0110000" when "0011",
		"0011001" when "0100",
		"0010010" when "0101",
		"0000010" when "0110",
		"1111000" when "0111",
		"0000000" when "1000",
		"0011000" when "1001",
		"0000110" when others;

end LOGICA_SIETE_SEGMENTOS;
